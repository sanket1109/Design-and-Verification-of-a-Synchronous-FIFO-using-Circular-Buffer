// FILES.svh

// packages
`include "packages/types.sv"

// interfaces
`include "interfaces/rtl_if.sv"

// rtl
`include "rtl/fifo.sv"
`include "rtl/top_rtl.sv"

// dv
`include "dv/top_tb.svh"

//coverage
`include "coverages.sv"
